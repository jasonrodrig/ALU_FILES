`define DATA_WIDTH 8
`define CMD_WIDTH  4  
`define no_of_transaction 5
`define DW 8
`define CW 4
parameter RESULT_WIDTH = 2 * `DATA_WIDTH ;
